.subckt DADFF_56ps D CK n07 n17 Q QN n09 n23 VDD VSS
MN001 n01 D VSS VSS				NMOS_VTL 	W=0.090000U L=0.050000U
MN002 n02 n03 VSS VSS 			NMOS_VTL 	W=0.220000U L=0.050000U
MN003 VSS n07 n04 VSS 			NMOS_VTL 	W=0.090000U L=0.050000U
MN004 n05 n02 n04 VSS 			NMOS_VTL 	W=0.090000U L=0.050000U
MN005 n06 n03 n05 VSS 			NMOS_VTL 	W=0.280000U L=0.050000U
MN006 n06 n01 VSS VSS 			NMOS_VTL 	W=0.280000U L=0.050000U
MN007 n07 n05 VSS VSS 			NMOS_VTL 	W=0.220000U L=0.050000U
MN008 VSS CK n03 VSS 			NMOS_VTL 	W=0.220000U L=0.050000U
MN009 n08 n05 VSS VSS 			NMOS_VTL 	W=0.220000U L=0.050000U
MN010 n09 n02 n08 VSS 			NMOS_VTL 	W=0.220000U L=0.050000U
MN011 n09 n03 n18 VSS 			NMOS_VTL 	W=0.090000U L=0.050000U
MN012 n18 n10 VSS VSS 			NMOS_VTL 	W=0.090000U L=0.050000U
MN013 VSS n09 n10 VSS 			NMOS_VTL 	W=0.220000U L=0.050000U
MN014 n15 n16 VSS VSS   		NMOS_VTL    W=0.220000U L=0.050000U
MN015 VSS n17 n21 VSS   		NMOS_VTL    W=0.090000U L=0.050000U
MN016 n20 n15 n21 VSS   		NMOS_VTL    W=0.090000U L=0.050000U
MN017 n19 n16 n20 VSS  			NMOS_VTL    W=0.280000U L=0.050000U
MN018 n24 Vref2 VSS VSS 		NMOS_VTL    W=0.210000U L=0.050000U
MN019 n19 n01 n24 VSS   		NMOS_VTL    W=0.280000U L=0.050000U
MN020 n17 n20 VSS VSS   		NMOS_VTL    W=0.220000U L=0.050000U
MN021 VSS CK n16 VSS    		NMOS_VTL    W=0.220000U L=0.050000U
MN022 n22 n20 VSS VSS   		NMOS_VTL    W=0.220000U L=0.050000U
MN023 n23 n15 n22 VSS  			NMOS_VTL    W=0.220000U L=0.050000U
MN024 n23 n16 n30 VSS 			NMOS_VTL    W=0.090000U L=0.050000U
MN025 n30 n29 VSS VSS  			NMOS_VTL    W=0.090000U L=0.050000U
MN026 VSS n23 n29 VSS  			NMOS_VTL    W=0.220000U L=0.050000U
MN027 n33 n23 n34 VSS   		NMOS_VTL 	W=0.210000U L=0.050000U
MN028 n34 n09 VSS VSS   		NMOS_VTL 	W=0.210000U L=0.050000U
MN029 QN n33 VSS VSS    		NMOS_VTL 	W=0.415000U L=0.050000U
MN030 Q QN VSS VSS      		NMOS_VTL 	W=0.415000U L=0.050000U
MN031 VSS Vref2 VSS VSS 		NMOS_VTL 	W=0.630000U L=0.050000U
MN032 VSS Vref4 VSS VSS 		NMOS_VTL 	W=0.630000U L=0.050000U
MP001 n33 n23 n32 VDD   		PMOS_VTL 	W=0.315000U L=0.050000U
MP002 n28 n29 VDD VDD 			PMOS_VTL    W=0.090000U L=0.050000U
MP003 VDD n23 n29 VDD  			PMOS_VTL    W=0.320000U L=0.050000U
MP004 n32 n09 VDD VDD   		PMOS_VTL 	W=0.315000U L=0.050000U
MP005 Q QN VDD VDD      		PMOS_VTL 	W=0.630000U L=0.050000U
MP006 QN n33 VDD VDD    		PMOS_VTL 	W=0.630000U L=0.050000U
MP007 n02 n03 VDD VDD 			PMOS_VTL 	W=0.320000U L=0.050000U
MP008 VDD n07 n11 VDD 			PMOS_VTL 	W=0.090000U L=0.050000U
MP009 n11 n03 n05 VDD 			PMOS_VTL 	W=0.090000U L=0.050000U
MP010 n05 n02 n12 VDD 			PMOS_VTL 	W=0.430000U L=0.050000U
MP011 n12 n01 VDD VDD 			PMOS_VTL 	W=0.430000U L=0.050000U
MP012 n07 n05 VDD VDD 			PMOS_VTL 	W=0.320000U L=0.050000U
MP013 VDD CK n03 VDD 			PMOS_VTL 	W=0.320000U L=0.050000U
MP014 n13 n05 VDD VDD 			PMOS_VTL 	W=0.320000U L=0.050000U
MP015 n09 n03 n13 VDD 			PMOS_VTL 	W=0.320000U L=0.050000U
MP016 n09 n02 n14 VDD 			PMOS_VTL 	W=0.090000U L=0.050000U
MP017 n01 D VDD VDD 			PMOS_VTL 	W=0.135000U L=0.050000U
MP018 n14 n10 VDD VDD 			PMOS_VTL 	W=0.090000U L=0.050000U
MP019 VDD n09 n10 VDD 			PMOS_VTL 	W=0.320000U L=0.050000U
MP020 n15 n16 VDD VDD   		PMOS_VTL    W=0.320000U L=0.050000U
MP021 VDD n17 n26 VDD   		PMOS_VTL    W=0.090000U L=0.050000U
MP022 n26 n16 n20 VDD  			PMOS_VTL    W=0.090000U L=0.050000U
MP023 n20 n15 n25 VDD   		PMOS_VTL    W=0.430000U L=0.050000U
MP024 n31 Vref4 VDD VDD 		PMOS_VTL    W=0.195000U L=0.050000U
MP025 n25 n01 n31 VDD   		PMOS_VTL    W=0.430000U L=0.050000U
MP026 n17 n20 VDD VDD   		PMOS_VTL    W=0.320000U L=0.050000U
MP027 VDD CK n16 VDD    		PMOS_VTL    W=0.320000U L=0.050000U
MP028 n27 n20 VDD VDD   		PMOS_VTL    W=0.320000U L=0.050000U
MP029 n23 n16 n27 VDD  			PMOS_VTL    W=0.320000U L=0.050000U
MP030 n23 n15 n28 VDD 			PMOS_VTL    W=0.090000U L=0.050000U
Mref00 VDD VDD Vref1 VSS		NMOS_VTL 	W=0.900000U L=0.050000U
Mref01 Vref1 Vref1 Vref2 VSS   	NMOS_VTL 	W=0.590000U L=0.050000U
Mref02 Vref2 Vref2 Vref3 VSS   	NMOS_VTL 	W=0.885000U L=0.050000U
Mref03 Vref3 Vref3 Vref4 VSS   	NMOS_VTL 	W=0.825000U L=0.050000U
Mref04 Vref4 Vref4 Vref5 VSS   	NMOS_VTL 	W=0.215000U L=0.050000U
Mref05 Vref5 Vref5 VSS VSS     	NMOS_VTL 	W=0.900000U L=0.050000U
.ends
